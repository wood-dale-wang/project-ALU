module ADD_32(
    input wire cin,
    input wire [31:0] a,
    input wire [31:0] b,
    output wire [31:0] res,
    output wire cout
  );

  wire [31:0] G;
  wire [31:0] P;
  wire [30:0] C;

  genvar i;

  generate
    for (i = 0; i < 32; i = i + 1)
    begin : add_bit
      and u_g_and(G[i],a[i],b[i]);
      or u_p_or(P[i],a[i],b[i]);
    end
  endgenerate

  // 产生cin相关位
  wire PxCIN[31:0];
  and u_and_p0cin(PxCIN[0],P[0],cin);
  and u_and_p1cin(PxCIN[1],P[1],P[0],cin);
  and u_and_p2cin(PxCIN[2],P[2],P[1],P[0],cin);
  and u_and_p3cin(PxCIN[3],P[3],P[2],P[1],P[0],cin);
  and u_and_p4cin(PxCIN[4],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p5cin(PxCIN[5],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p6cin(PxCIN[6],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p7cin(PxCIN[7],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p8cin(PxCIN[8],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p9cin(PxCIN[9],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p10cin(PxCIN[10],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p11cin(PxCIN[11],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p12cin(PxCIN[12],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p13cin(PxCIN[13],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p14cin(PxCIN[14],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p15cin(PxCIN[15],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p16cin(PxCIN[16],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p17cin(PxCIN[17],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p18cin(PxCIN[18],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p19cin(PxCIN[19],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p20cin(PxCIN[20],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p21cin(PxCIN[21],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p22cin(PxCIN[22],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p23cin(PxCIN[23],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p24cin(PxCIN[24],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p25cin(PxCIN[25],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p26cin(PxCIN[26],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p27cin(PxCIN[27],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p28cin(PxCIN[28],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p29cin(PxCIN[29],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p30cin(PxCIN[30],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);
  and u_and_p31cin(PxCIN[31],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0],cin);


  // 产生G0相关位
  wire PxG0[30:0];
  and u_and_p1g0(PxG0[0],P[1],G[0]);
  and u_and_p2g0(PxG0[1],P[2],P[1],G[0]);
  and u_and_p3g0(PxG0[2],P[3],P[2],P[1],G[0]);
  and u_and_p4g0(PxG0[3],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p5g0(PxG0[4],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p6g0(PxG0[5],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p7g0(PxG0[6],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p8g0(PxG0[7],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p9g0(PxG0[8],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p10g0(PxG0[9],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p11g0(PxG0[10],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p12g0(PxG0[11],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p13g0(PxG0[12],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p14g0(PxG0[13],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p15g0(PxG0[14],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p16g0(PxG0[15],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p17g0(PxG0[16],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p18g0(PxG0[17],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p19g0(PxG0[18],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p20g0(PxG0[19],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p21g0(PxG0[20],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p22g0(PxG0[21],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p23g0(PxG0[22],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p24g0(PxG0[23],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p25g0(PxG0[24],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p26g0(PxG0[25],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p27g0(PxG0[26],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p28g0(PxG0[27],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p29g0(PxG0[28],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p30g0(PxG0[29],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  and u_and_p31g0(PxG0[30],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],P[1],G[0]);
  wire PxG1[29:0];
  and u_and_p2g1(PxG1[0],P[2],G[1]);
  and u_and_p3g1(PxG1[1],P[3],P[2],G[1]);
  and u_and_p4g1(PxG1[2],P[4],P[3],P[2],G[1]);
  and u_and_p5g1(PxG1[3],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p6g1(PxG1[4],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p7g1(PxG1[5],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p8g1(PxG1[6],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p9g1(PxG1[7],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p10g1(PxG1[8],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p11g1(PxG1[9],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p12g1(PxG1[10],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p13g1(PxG1[11],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p14g1(PxG1[12],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p15g1(PxG1[13],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p16g1(PxG1[14],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p17g1(PxG1[15],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p18g1(PxG1[16],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p19g1(PxG1[17],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p20g1(PxG1[18],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p21g1(PxG1[19],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p22g1(PxG1[20],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p23g1(PxG1[21],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p24g1(PxG1[22],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p25g1(PxG1[23],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p26g1(PxG1[24],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p27g1(PxG1[25],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p28g1(PxG1[26],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p29g1(PxG1[27],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p30g1(PxG1[28],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  and u_and_p31g1(PxG1[29],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],P[2],G[1]);
  wire PxG2[28:0];
  and u_and_p3g2(PxG2[0],P[3],G[2]);
  and u_and_p4g2(PxG2[1],P[4],P[3],G[2]);
  and u_and_p5g2(PxG2[2],P[5],P[4],P[3],G[2]);
  and u_and_p6g2(PxG2[3],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p7g2(PxG2[4],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p8g2(PxG2[5],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p9g2(PxG2[6],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p10g2(PxG2[7],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p11g2(PxG2[8],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p12g2(PxG2[9],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p13g2(PxG2[10],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p14g2(PxG2[11],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p15g2(PxG2[12],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p16g2(PxG2[13],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p17g2(PxG2[14],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p18g2(PxG2[15],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p19g2(PxG2[16],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p20g2(PxG2[17],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p21g2(PxG2[18],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p22g2(PxG2[19],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p23g2(PxG2[20],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p24g2(PxG2[21],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p25g2(PxG2[22],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p26g2(PxG2[23],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p27g2(PxG2[24],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p28g2(PxG2[25],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p29g2(PxG2[26],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p30g2(PxG2[27],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  and u_and_p31g2(PxG2[28],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],P[3],G[2]);
  wire PxG3[27:0];
  and u_and_p4g3(PxG3[0],P[4],G[3]);
  and u_and_p5g3(PxG3[1],P[5],P[4],G[3]);
  and u_and_p6g3(PxG3[2],P[6],P[5],P[4],G[3]);
  and u_and_p7g3(PxG3[3],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p8g3(PxG3[4],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p9g3(PxG3[5],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p10g3(PxG3[6],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p11g3(PxG3[7],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p12g3(PxG3[8],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p13g3(PxG3[9],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p14g3(PxG3[10],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p15g3(PxG3[11],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p16g3(PxG3[12],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p17g3(PxG3[13],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p18g3(PxG3[14],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p19g3(PxG3[15],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p20g3(PxG3[16],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p21g3(PxG3[17],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p22g3(PxG3[18],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p23g3(PxG3[19],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p24g3(PxG3[20],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p25g3(PxG3[21],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p26g3(PxG3[22],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p27g3(PxG3[23],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p28g3(PxG3[24],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p29g3(PxG3[25],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p30g3(PxG3[26],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  and u_and_p31g3(PxG3[27],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],P[4],G[3]);
  wire PxG4[26:0];
  and u_and_p5g4(PxG4[0],P[5],G[4]);
  and u_and_p6g4(PxG4[1],P[6],P[5],G[4]);
  and u_and_p7g4(PxG4[2],P[7],P[6],P[5],G[4]);
  and u_and_p8g4(PxG4[3],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p9g4(PxG4[4],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p10g4(PxG4[5],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p11g4(PxG4[6],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p12g4(PxG4[7],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p13g4(PxG4[8],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p14g4(PxG4[9],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p15g4(PxG4[10],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p16g4(PxG4[11],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p17g4(PxG4[12],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p18g4(PxG4[13],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p19g4(PxG4[14],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p20g4(PxG4[15],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p21g4(PxG4[16],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p22g4(PxG4[17],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p23g4(PxG4[18],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p24g4(PxG4[19],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p25g4(PxG4[20],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p26g4(PxG4[21],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p27g4(PxG4[22],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p28g4(PxG4[23],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p29g4(PxG4[24],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p30g4(PxG4[25],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  and u_and_p31g4(PxG4[26],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],P[5],G[4]);
  wire PxG5[25:0];
  and u_and_p6g5(PxG5[0],P[6],G[5]);
  and u_and_p7g5(PxG5[1],P[7],P[6],G[5]);
  and u_and_p8g5(PxG5[2],P[8],P[7],P[6],G[5]);
  and u_and_p9g5(PxG5[3],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p10g5(PxG5[4],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p11g5(PxG5[5],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p12g5(PxG5[6],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p13g5(PxG5[7],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p14g5(PxG5[8],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p15g5(PxG5[9],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p16g5(PxG5[10],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p17g5(PxG5[11],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p18g5(PxG5[12],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p19g5(PxG5[13],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p20g5(PxG5[14],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p21g5(PxG5[15],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p22g5(PxG5[16],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p23g5(PxG5[17],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p24g5(PxG5[18],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p25g5(PxG5[19],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p26g5(PxG5[20],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p27g5(PxG5[21],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p28g5(PxG5[22],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p29g5(PxG5[23],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p30g5(PxG5[24],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  and u_and_p31g5(PxG5[25],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],P[6],G[5]);
  wire PxG6[24:0];
  and u_and_p7g6(PxG6[0],P[7],G[6]);
  and u_and_p8g6(PxG6[1],P[8],P[7],G[6]);
  and u_and_p9g6(PxG6[2],P[9],P[8],P[7],G[6]);
  and u_and_p10g6(PxG6[3],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p11g6(PxG6[4],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p12g6(PxG6[5],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p13g6(PxG6[6],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p14g6(PxG6[7],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p15g6(PxG6[8],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p16g6(PxG6[9],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p17g6(PxG6[10],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p18g6(PxG6[11],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p19g6(PxG6[12],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p20g6(PxG6[13],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p21g6(PxG6[14],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p22g6(PxG6[15],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p23g6(PxG6[16],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p24g6(PxG6[17],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p25g6(PxG6[18],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p26g6(PxG6[19],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p27g6(PxG6[20],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p28g6(PxG6[21],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p29g6(PxG6[22],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p30g6(PxG6[23],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  and u_and_p31g6(PxG6[24],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],P[7],G[6]);
  wire PxG7[23:0];
  and u_and_p8g7(PxG7[0],P[8],G[7]);
  and u_and_p9g7(PxG7[1],P[9],P[8],G[7]);
  and u_and_p10g7(PxG7[2],P[10],P[9],P[8],G[7]);
  and u_and_p11g7(PxG7[3],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p12g7(PxG7[4],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p13g7(PxG7[5],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p14g7(PxG7[6],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p15g7(PxG7[7],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p16g7(PxG7[8],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p17g7(PxG7[9],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p18g7(PxG7[10],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p19g7(PxG7[11],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p20g7(PxG7[12],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p21g7(PxG7[13],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p22g7(PxG7[14],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p23g7(PxG7[15],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p24g7(PxG7[16],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p25g7(PxG7[17],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p26g7(PxG7[18],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p27g7(PxG7[19],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p28g7(PxG7[20],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p29g7(PxG7[21],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p30g7(PxG7[22],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  and u_and_p31g7(PxG7[23],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],P[8],G[7]);
  wire PxG8[22:0];
  and u_and_p9g8(PxG8[0],P[9],G[8]);
  and u_and_p10g8(PxG8[1],P[10],P[9],G[8]);
  and u_and_p11g8(PxG8[2],P[11],P[10],P[9],G[8]);
  and u_and_p12g8(PxG8[3],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p13g8(PxG8[4],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p14g8(PxG8[5],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p15g8(PxG8[6],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p16g8(PxG8[7],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p17g8(PxG8[8],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p18g8(PxG8[9],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p19g8(PxG8[10],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p20g8(PxG8[11],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p21g8(PxG8[12],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p22g8(PxG8[13],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p23g8(PxG8[14],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p24g8(PxG8[15],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p25g8(PxG8[16],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p26g8(PxG8[17],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p27g8(PxG8[18],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p28g8(PxG8[19],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p29g8(PxG8[20],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p30g8(PxG8[21],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  and u_and_p31g8(PxG8[22],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],P[9],G[8]);
  wire PxG9[21:0];
  and u_and_p10g9(PxG9[0],P[10],G[9]);
  and u_and_p11g9(PxG9[1],P[11],P[10],G[9]);
  and u_and_p12g9(PxG9[2],P[12],P[11],P[10],G[9]);
  and u_and_p13g9(PxG9[3],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p14g9(PxG9[4],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p15g9(PxG9[5],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p16g9(PxG9[6],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p17g9(PxG9[7],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p18g9(PxG9[8],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p19g9(PxG9[9],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p20g9(PxG9[10],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p21g9(PxG9[11],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p22g9(PxG9[12],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p23g9(PxG9[13],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p24g9(PxG9[14],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p25g9(PxG9[15],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p26g9(PxG9[16],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p27g9(PxG9[17],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p28g9(PxG9[18],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p29g9(PxG9[19],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p30g9(PxG9[20],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  and u_and_p31g9(PxG9[21],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],P[10],G[9]);
  wire PxG10[20:0];
  and u_and_p11g10(PxG10[0],P[11],G[10]);
  and u_and_p12g10(PxG10[1],P[12],P[11],G[10]);
  and u_and_p13g10(PxG10[2],P[13],P[12],P[11],G[10]);
  and u_and_p14g10(PxG10[3],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p15g10(PxG10[4],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p16g10(PxG10[5],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p17g10(PxG10[6],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p18g10(PxG10[7],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p19g10(PxG10[8],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p20g10(PxG10[9],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p21g10(PxG10[10],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p22g10(PxG10[11],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p23g10(PxG10[12],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p24g10(PxG10[13],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p25g10(PxG10[14],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p26g10(PxG10[15],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p27g10(PxG10[16],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p28g10(PxG10[17],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p29g10(PxG10[18],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p30g10(PxG10[19],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  and u_and_p31g10(PxG10[20],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],P[11],G[10]);
  wire PxG11[19:0];
  and u_and_p12g11(PxG11[0],P[12],G[11]);
  and u_and_p13g11(PxG11[1],P[13],P[12],G[11]);
  and u_and_p14g11(PxG11[2],P[14],P[13],P[12],G[11]);
  and u_and_p15g11(PxG11[3],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p16g11(PxG11[4],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p17g11(PxG11[5],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p18g11(PxG11[6],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p19g11(PxG11[7],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p20g11(PxG11[8],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p21g11(PxG11[9],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p22g11(PxG11[10],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p23g11(PxG11[11],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p24g11(PxG11[12],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p25g11(PxG11[13],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p26g11(PxG11[14],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p27g11(PxG11[15],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p28g11(PxG11[16],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p29g11(PxG11[17],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p30g11(PxG11[18],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  and u_and_p31g11(PxG11[19],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],P[12],G[11]);
  wire PxG12[18:0];
  and u_and_p13g12(PxG12[0],P[13],G[12]);
  and u_and_p14g12(PxG12[1],P[14],P[13],G[12]);
  and u_and_p15g12(PxG12[2],P[15],P[14],P[13],G[12]);
  and u_and_p16g12(PxG12[3],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p17g12(PxG12[4],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p18g12(PxG12[5],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p19g12(PxG12[6],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p20g12(PxG12[7],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p21g12(PxG12[8],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p22g12(PxG12[9],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p23g12(PxG12[10],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p24g12(PxG12[11],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p25g12(PxG12[12],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p26g12(PxG12[13],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p27g12(PxG12[14],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p28g12(PxG12[15],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p29g12(PxG12[16],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p30g12(PxG12[17],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  and u_and_p31g12(PxG12[18],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],P[13],G[12]);
  wire PxG13[17:0];
  and u_and_p14g13(PxG13[0],P[14],G[13]);
  and u_and_p15g13(PxG13[1],P[15],P[14],G[13]);
  and u_and_p16g13(PxG13[2],P[16],P[15],P[14],G[13]);
  and u_and_p17g13(PxG13[3],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p18g13(PxG13[4],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p19g13(PxG13[5],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p20g13(PxG13[6],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p21g13(PxG13[7],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p22g13(PxG13[8],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p23g13(PxG13[9],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p24g13(PxG13[10],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p25g13(PxG13[11],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p26g13(PxG13[12],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p27g13(PxG13[13],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p28g13(PxG13[14],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p29g13(PxG13[15],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p30g13(PxG13[16],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  and u_and_p31g13(PxG13[17],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],P[14],G[13]);
  wire PxG14[16:0];
  and u_and_p15g14(PxG14[0],P[15],G[14]);
  and u_and_p16g14(PxG14[1],P[16],P[15],G[14]);
  and u_and_p17g14(PxG14[2],P[17],P[16],P[15],G[14]);
  and u_and_p18g14(PxG14[3],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p19g14(PxG14[4],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p20g14(PxG14[5],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p21g14(PxG14[6],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p22g14(PxG14[7],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p23g14(PxG14[8],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p24g14(PxG14[9],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p25g14(PxG14[10],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p26g14(PxG14[11],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p27g14(PxG14[12],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p28g14(PxG14[13],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p29g14(PxG14[14],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p30g14(PxG14[15],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  and u_and_p31g14(PxG14[16],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],P[15],G[14]);
  wire PxG15[15:0];
  and u_and_p16g15(PxG15[0],P[16],G[15]);
  and u_and_p17g15(PxG15[1],P[17],P[16],G[15]);
  and u_and_p18g15(PxG15[2],P[18],P[17],P[16],G[15]);
  and u_and_p19g15(PxG15[3],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p20g15(PxG15[4],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p21g15(PxG15[5],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p22g15(PxG15[6],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p23g15(PxG15[7],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p24g15(PxG15[8],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p25g15(PxG15[9],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p26g15(PxG15[10],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p27g15(PxG15[11],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p28g15(PxG15[12],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p29g15(PxG15[13],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p30g15(PxG15[14],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  and u_and_p31g15(PxG15[15],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],P[16],G[15]);
  wire PxG16[14:0];
  and u_and_p17g16(PxG16[0],P[17],G[16]);
  and u_and_p18g16(PxG16[1],P[18],P[17],G[16]);
  and u_and_p19g16(PxG16[2],P[19],P[18],P[17],G[16]);
  and u_and_p20g16(PxG16[3],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p21g16(PxG16[4],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p22g16(PxG16[5],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p23g16(PxG16[6],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p24g16(PxG16[7],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p25g16(PxG16[8],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p26g16(PxG16[9],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p27g16(PxG16[10],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p28g16(PxG16[11],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p29g16(PxG16[12],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p30g16(PxG16[13],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  and u_and_p31g16(PxG16[14],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],P[17],G[16]);
  wire PxG17[13:0];
  and u_and_p18g17(PxG17[0],P[18],G[17]);
  and u_and_p19g17(PxG17[1],P[19],P[18],G[17]);
  and u_and_p20g17(PxG17[2],P[20],P[19],P[18],G[17]);
  and u_and_p21g17(PxG17[3],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p22g17(PxG17[4],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p23g17(PxG17[5],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p24g17(PxG17[6],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p25g17(PxG17[7],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p26g17(PxG17[8],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p27g17(PxG17[9],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p28g17(PxG17[10],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p29g17(PxG17[11],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p30g17(PxG17[12],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  and u_and_p31g17(PxG17[13],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],P[18],G[17]);
  wire PxG18[12:0];
  and u_and_p19g18(PxG18[0],P[19],G[18]);
  and u_and_p20g18(PxG18[1],P[20],P[19],G[18]);
  and u_and_p21g18(PxG18[2],P[21],P[20],P[19],G[18]);
  and u_and_p22g18(PxG18[3],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p23g18(PxG18[4],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p24g18(PxG18[5],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p25g18(PxG18[6],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p26g18(PxG18[7],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p27g18(PxG18[8],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p28g18(PxG18[9],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p29g18(PxG18[10],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p30g18(PxG18[11],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  and u_and_p31g18(PxG18[12],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],P[19],G[18]);
  wire PxG19[11:0];
  and u_and_p20g19(PxG19[0],P[20],G[19]);
  and u_and_p21g19(PxG19[1],P[21],P[20],G[19]);
  and u_and_p22g19(PxG19[2],P[22],P[21],P[20],G[19]);
  and u_and_p23g19(PxG19[3],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p24g19(PxG19[4],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p25g19(PxG19[5],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p26g19(PxG19[6],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p27g19(PxG19[7],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p28g19(PxG19[8],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p29g19(PxG19[9],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p30g19(PxG19[10],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  and u_and_p31g19(PxG19[11],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],P[20],G[19]);
  wire PxG20[10:0];
  and u_and_p21g20(PxG20[0],P[21],G[20]);
  and u_and_p22g20(PxG20[1],P[22],P[21],G[20]);
  and u_and_p23g20(PxG20[2],P[23],P[22],P[21],G[20]);
  and u_and_p24g20(PxG20[3],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p25g20(PxG20[4],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p26g20(PxG20[5],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p27g20(PxG20[6],P[27],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p28g20(PxG20[7],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p29g20(PxG20[8],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p30g20(PxG20[9],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  and u_and_p31g20(PxG20[10],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],P[21],G[20]);
  wire PxG21[9:0];
  and u_and_p22g21(PxG21[0],P[22],G[21]);
  and u_and_p23g21(PxG21[1],P[23],P[22],G[21]);
  and u_and_p24g21(PxG21[2],P[24],P[23],P[22],G[21]);
  and u_and_p25g21(PxG21[3],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p26g21(PxG21[4],P[26],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p27g21(PxG21[5],P[27],P[26],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p28g21(PxG21[6],P[28],P[27],P[26],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p29g21(PxG21[7],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p30g21(PxG21[8],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],G[21]);
  and u_and_p31g21(PxG21[9],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],P[22],G[21]);
  wire PxG22[8:0];
  and u_and_p23g22(PxG22[0],P[23],G[22]);
  and u_and_p24g22(PxG22[1],P[24],P[23],G[22]);
  and u_and_p25g22(PxG22[2],P[25],P[24],P[23],G[22]);
  and u_and_p26g22(PxG22[3],P[26],P[25],P[24],P[23],G[22]);
  and u_and_p27g22(PxG22[4],P[27],P[26],P[25],P[24],P[23],G[22]);
  and u_and_p28g22(PxG22[5],P[28],P[27],P[26],P[25],P[24],P[23],G[22]);
  and u_and_p29g22(PxG22[6],P[29],P[28],P[27],P[26],P[25],P[24],P[23],G[22]);
  and u_and_p30g22(PxG22[7],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],G[22]);
  and u_and_p31g22(PxG22[8],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],P[23],G[22]);
  wire PxG23[7:0];
  and u_and_p24g23(PxG23[0],P[24],G[23]);
  and u_and_p25g23(PxG23[1],P[25],P[24],G[23]);
  and u_and_p26g23(PxG23[2],P[26],P[25],P[24],G[23]);
  and u_and_p27g23(PxG23[3],P[27],P[26],P[25],P[24],G[23]);
  and u_and_p28g23(PxG23[4],P[28],P[27],P[26],P[25],P[24],G[23]);
  and u_and_p29g23(PxG23[5],P[29],P[28],P[27],P[26],P[25],P[24],G[23]);
  and u_and_p30g23(PxG23[6],P[30],P[29],P[28],P[27],P[26],P[25],P[24],G[23]);
  and u_and_p31g23(PxG23[7],P[31],P[30],P[29],P[28],P[27],P[26],P[25],P[24],G[23]);
  wire PxG24[6:0];
  and u_and_p25g24(PxG24[0],P[25],G[24]);
  and u_and_p26g24(PxG24[1],P[26],P[25],G[24]);
  and u_and_p27g24(PxG24[2],P[27],P[26],P[25],G[24]);
  and u_and_p28g24(PxG24[3],P[28],P[27],P[26],P[25],G[24]);
  and u_and_p29g24(PxG24[4],P[29],P[28],P[27],P[26],P[25],G[24]);
  and u_and_p30g24(PxG24[5],P[30],P[29],P[28],P[27],P[26],P[25],G[24]);
  and u_and_p31g24(PxG24[6],P[31],P[30],P[29],P[28],P[27],P[26],P[25],G[24]);
  wire PxG25[5:0];
  and u_and_p26g25(PxG25[0],P[26],G[25]);
  and u_and_p27g25(PxG25[1],P[27],P[26],G[25]);
  and u_and_p28g25(PxG25[2],P[28],P[27],P[26],G[25]);
  and u_and_p29g25(PxG25[3],P[29],P[28],P[27],P[26],G[25]);
  and u_and_p30g25(PxG25[4],P[30],P[29],P[28],P[27],P[26],G[25]);
  and u_and_p31g25(PxG25[5],P[31],P[30],P[29],P[28],P[27],P[26],G[25]);
  wire PxG26[4:0];
  and u_and_p27g26(PxG26[0],P[27],G[26]);
  and u_and_p28g26(PxG26[1],P[28],P[27],G[26]);
  and u_and_p29g26(PxG26[2],P[29],P[28],P[27],G[26]);
  and u_and_p30g26(PxG26[3],P[30],P[29],P[28],P[27],G[26]);
  and u_and_p31g26(PxG26[4],P[31],P[30],P[29],P[28],P[27],G[26]);
  wire PxG27[3:0];
  and u_and_p28g27(PxG27[0],P[28],G[27]);
  and u_and_p29g27(PxG27[1],P[29],P[28],G[27]);
  and u_and_p30g27(PxG27[2],P[30],P[29],P[28],G[27]);
  and u_and_p31g27(PxG27[3],P[31],P[30],P[29],P[28],G[27]);
  wire PxG28[2:0];
  and u_and_p29g28(PxG28[0],P[29],G[28]);
  and u_and_p30g28(PxG28[1],P[30],P[29],G[28]);
  and u_and_p31g28(PxG28[2],P[31],P[30],P[29],G[28]);
  wire PxG29[1:0];
  and u_and_p30g29(PxG29[0],P[30],G[29]);
  and u_and_p31g29(PxG29[1],P[31],P[30],G[29]);
  wire PxG30;
  and u_and_p31g30(PxG30,P[31],G[30]);

  // 产生C
  or u_or_c0(C[0],G[0],PxCIN[0]);
  or u_or_c1(C[1],G[1],PxG0[0],PxCIN[1]);
  or u_or_c2(C[2],G[2],PxG1[0],PxG0[1],PxCIN[2]);
  or u_or_c3(C[3],G[3],PxG2[0],PxG1[1],PxG0[2],PxCIN[3]);
  or u_or_c4(C[4],G[4],PxG3[0],PxG2[1],PxG1[2],PxG0[3],PxCIN[4]);
  or u_or_c5(C[5],G[5],PxG4[0],PxG3[1],PxG2[2],PxG1[3],PxG0[4],PxCIN[5]);
  or u_or_c6(C[6],G[6],PxG5[0],PxG4[1],PxG3[2],PxG2[3],PxG1[4],PxG0[5],PxCIN[6]);
  or u_or_c7(C[7],G[7],PxG6[0],PxG5[1],PxG4[2],PxG3[3],PxG2[4],PxG1[5],PxG0[6],PxCIN[7]);
  or u_or_c8(C[8],G[8],PxG7[0],PxG6[1],PxG5[2],PxG4[3],PxG3[4],PxG2[5],PxG1[6],PxG0[7],PxCIN[8]);
  or u_or_c9(C[9],G[9],PxG8[0],PxG7[1],PxG6[2],PxG5[3],PxG4[4],PxG3[5],PxG2[6],PxG1[7],PxG0[8],PxCIN[9]);
  or u_or_c10(C[10],G[10],PxG9[0],PxG8[1],PxG7[2],PxG6[3],PxG5[4],PxG4[5],PxG3[6],PxG2[7],PxG1[8],PxG0[9],PxCIN[10]);
  or u_or_c11(C[11],G[11],PxG10[0],PxG9[1],PxG8[2],PxG7[3],PxG6[4],PxG5[5],PxG4[6],PxG3[7],PxG2[8],PxG1[9],PxG0[10],PxCIN[11]);
  or u_or_c12(C[12],G[12],PxG11[0],PxG10[1],PxG9[2],PxG8[3],PxG7[4],PxG6[5],PxG5[6],PxG4[7],PxG3[8],PxG2[9],PxG1[10],PxG0[11],PxCIN[12]);
  or u_or_c13(C[13],G[13],PxG12[0],PxG11[1],PxG10[2],PxG9[3],PxG8[4],PxG7[5],PxG6[6],PxG5[7],PxG4[8],PxG3[9],PxG2[10],PxG1[11],PxG0[12],PxCIN[13]);
  or u_or_c14(C[14],G[14],PxG13[0],PxG12[1],PxG11[2],PxG10[3],PxG9[4],PxG8[5],PxG7[6],PxG6[7],PxG5[8],PxG4[9],PxG3[10],PxG2[11],PxG1[12],PxG0[13],PxCIN[14]);
  or u_or_c15(C[15],G[15],PxG14[0],PxG13[1],PxG12[2],PxG11[3],PxG10[4],PxG9[5],PxG8[6],PxG7[7],PxG6[8],PxG5[9],PxG4[10],PxG3[11],PxG2[12],PxG1[13],PxG0[14],PxCIN[15]);
  or u_or_c16(C[16],G[16],PxG15[0],PxG14[1],PxG13[2],PxG12[3],PxG11[4],PxG10[5],PxG9[6],PxG8[7],PxG7[8],PxG6[9],PxG5[10],PxG4[11],PxG3[12],PxG2[13],PxG1[14],PxG0[15],PxCIN[16]);
  or u_or_c17(C[17],G[17],PxG16[0],PxG15[1],PxG14[2],PxG13[3],PxG12[4],PxG11[5],PxG10[6],PxG9[7],PxG8[8],PxG7[9],PxG6[10],PxG5[11],PxG4[12],PxG3[13],PxG2[14],PxG1[15],PxG0[16],PxCIN[17]);
  or u_or_c18(C[18],G[18],PxG17[0],PxG16[1],PxG15[2],PxG14[3],PxG13[4],PxG12[5],PxG11[6],PxG10[7],PxG9[8],PxG8[9],PxG7[10],PxG6[11],PxG5[12],PxG4[13],PxG3[14],PxG2[15],PxG1[16],PxG0[17],PxCIN[18]);
  or u_or_c19(C[19],G[19],PxG18[0],PxG17[1],PxG16[2],PxG15[3],PxG14[4],PxG13[5],PxG12[6],PxG11[7],PxG10[8],PxG9[9],PxG8[10],PxG7[11],PxG6[12],PxG5[13],PxG4[14],PxG3[15],PxG2[16],PxG1[17],PxG0[18],PxCIN[19]);
  or u_or_c20(C[20],G[20],PxG19[0],PxG18[1],PxG17[2],PxG16[3],PxG15[4],PxG14[5],PxG13[6],PxG12[7],PxG11[8],PxG10[9],PxG9[10],PxG8[11],PxG7[12],PxG6[13],PxG5[14],PxG4[15],PxG3[16],PxG2[17],PxG1[18],PxG0[19],PxCIN[20]);
  or u_or_c21(C[21],G[21],PxG20[0],PxG19[1],PxG18[2],PxG17[3],PxG16[4],PxG15[5],PxG14[6],PxG13[7],PxG12[8],PxG11[9],PxG10[10],PxG9[11],PxG8[12],PxG7[13],PxG6[14],PxG5[15],PxG4[16],PxG3[17],PxG2[18],PxG1[19],PxG0[20],PxCIN[21]);
  or u_or_c22(C[22],G[22],PxG21[0],PxG20[1],PxG19[2],PxG18[3],PxG17[4],PxG16[5],PxG15[6],PxG14[7],PxG13[8],PxG12[9],PxG11[10],PxG10[11],PxG9[12],PxG8[13],PxG7[14],PxG6[15],PxG5[16],PxG4[17],PxG3[18],PxG2[19],PxG1[20],PxG0[21],PxCIN[22]);
  or u_or_c23(C[23],G[23],PxG22[0],PxG21[1],PxG20[2],PxG19[3],PxG18[4],PxG17[5],PxG16[6],PxG15[7],PxG14[8],PxG13[9],PxG12[10],PxG11[11],PxG10[12],PxG9[13],PxG8[14],PxG7[15],PxG6[16],PxG5[17],PxG4[18],PxG3[19],PxG2[20],PxG1[21],PxG0[22],PxCIN[23]);
  or u_or_c24(C[24],G[24],PxG23[0],PxG22[1],PxG21[2],PxG20[3],PxG19[4],PxG18[5],PxG17[6],PxG16[7],PxG15[8],PxG14[9],PxG13[10],PxG12[11],PxG11[12],PxG10[13],PxG9[14],PxG8[15],PxG7[16],PxG6[17],PxG5[18],PxG4[19],PxG3[20],PxG2[21],PxG1[22],PxG0[23],PxCIN[24]);
  or u_or_c25(C[25],G[25],PxG24[0],PxG23[1],PxG22[2],PxG21[3],PxG20[4],PxG19[5],PxG18[6],PxG17[7],PxG16[8],PxG15[9],PxG14[10],PxG13[11],PxG12[12],PxG11[13],PxG10[14],PxG9[15],PxG8[16],PxG7[17],PxG6[18],PxG5[19],PxG4[20],PxG3[21],PxG2[22],PxG1[23],PxG0[24],PxCIN[25]);
  or u_or_c26(C[26],G[26],PxG25[0],PxG24[1],PxG23[2],PxG22[3],PxG21[4],PxG20[5],PxG19[6],PxG18[7],PxG17[8],PxG16[9],PxG15[10],PxG14[11],PxG13[12],PxG12[13],PxG11[14],PxG10[15],PxG9[16],PxG8[17],PxG7[18],PxG6[19],PxG5[20],PxG4[21],PxG3[22],PxG2[23],PxG1[24],PxG0[25],PxCIN[26]);
  or u_or_c27(C[27],G[27],PxG26[0],PxG25[1],PxG24[2],PxG23[3],PxG22[4],PxG21[5],PxG20[6],PxG19[7],PxG18[8],PxG17[9],PxG16[10],PxG15[11],PxG14[12],PxG13[13],PxG12[14],PxG11[15],PxG10[16],PxG9[17],PxG8[18],PxG7[19],PxG6[20],PxG5[21],PxG4[22],PxG3[23],PxG2[24],PxG1[25],PxG0[26],PxCIN[27]);
  or u_or_c28(C[28],G[28],PxG27[0],PxG26[1],PxG25[2],PxG24[3],PxG23[4],PxG22[5],PxG21[6],PxG20[7],PxG19[8],PxG18[9],PxG17[10],PxG16[11],PxG15[12],PxG14[13],PxG13[14],PxG12[15],PxG11[16],PxG10[17],PxG9[18],PxG8[19],PxG7[20],PxG6[21],PxG5[22],PxG4[23],PxG3[24],PxG2[25],PxG1[26],PxG0[27],PxCIN[28]);
  or u_or_c29(C[29],G[29],PxG28[0],PxG27[1],PxG26[2],PxG25[3],PxG24[4],PxG23[5],PxG22[6],PxG21[7],PxG20[8],PxG19[9],PxG18[10],PxG17[11],PxG16[12],PxG15[13],PxG14[14],PxG13[15],PxG12[16],PxG11[17],PxG10[18],PxG9[19],PxG8[20],PxG7[21],PxG6[22],PxG5[23],PxG4[24],PxG3[25],PxG2[26],PxG1[27],PxG0[28],PxCIN[29]);
  or u_or_c30(C[30],G[30],PxG29[0],PxG28[1],PxG27[2],PxG26[3],PxG25[4],PxG24[5],PxG23[6],PxG22[7],PxG21[8],PxG20[9],PxG19[10],PxG18[11],PxG17[12],PxG16[13],PxG15[14],PxG14[15],PxG13[16],PxG12[17],PxG11[18],PxG10[19],PxG9[20],PxG8[21],PxG7[22],PxG6[23],PxG5[24],PxG4[25],PxG3[26],PxG2[27],PxG1[28],PxG0[29],PxCIN[30]);
  or u_or_c31(cout,G[31],PxG30,PxG29[1],PxG28[2],PxG27[3],PxG26[4],PxG25[5],PxG24[6],PxG23[7],PxG22[8],PxG21[9],PxG20[10],PxG19[11],PxG18[12],PxG17[13],PxG16[14],PxG15[15],PxG14[16],PxG13[17],PxG12[18],PxG11[19],PxG10[20],PxG9[21],PxG8[22],PxG7[23],PxG6[24],PxG5[25],PxG4[26],PxG3[27],PxG2[28],PxG1[29],PxG0[30],PxCIN[31]);

  // 产生res
  xor u_xor_r0(res[0],a[0],b[0],cin);
  xor u_xor_r1(res[1],a[1],b[1],C[0]);
  xor u_xor_r2(res[2],a[2],b[2],C[1]);
  xor u_xor_r3(res[3],a[3],b[3],C[2]);
  xor u_xor_r4(res[4],a[4],b[4],C[3]);
  xor u_xor_r5(res[5],a[5],b[5],C[4]);
  xor u_xor_r6(res[6],a[6],b[6],C[5]);
  xor u_xor_r7(res[7],a[7],b[7],C[6]);
  xor u_xor_r8(res[8],a[8],b[8],C[7]);
  xor u_xor_r9(res[9],a[9],b[9],C[8]);
  xor u_xor_r10(res[10],a[10],b[10],C[9]);
  xor u_xor_r11(res[11],a[11],b[11],C[10]);
  xor u_xor_r12(res[12],a[12],b[12],C[11]);
  xor u_xor_r13(res[13],a[13],b[13],C[12]);
  xor u_xor_r14(res[14],a[14],b[14],C[13]);
  xor u_xor_r15(res[15],a[15],b[15],C[14]);
  xor u_xor_r16(res[16],a[16],b[16],C[15]);
  xor u_xor_r17(res[17],a[17],b[17],C[16]);
  xor u_xor_r18(res[18],a[18],b[18],C[17]);
  xor u_xor_r19(res[19],a[19],b[19],C[18]);
  xor u_xor_r20(res[20],a[20],b[20],C[19]);
  xor u_xor_r21(res[21],a[21],b[21],C[20]);
  xor u_xor_r22(res[22],a[22],b[22],C[21]);
  xor u_xor_r23(res[23],a[23],b[23],C[22]);
  xor u_xor_r24(res[24],a[24],b[24],C[23]);
  xor u_xor_r25(res[25],a[25],b[25],C[24]);
  xor u_xor_r26(res[26],a[26],b[26],C[25]);
  xor u_xor_r27(res[27],a[27],b[27],C[26]);
  xor u_xor_r28(res[28],a[28],b[28],C[27]);
  xor u_xor_r29(res[29],a[29],b[29],C[28]);
  xor u_xor_r30(res[30],a[30],b[30],C[29]);
  xor u_xor_r31(res[31],a[31],b[31],C[30]);

endmodule
